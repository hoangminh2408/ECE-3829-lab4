`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/24/2019 05:15:00 PM
// Design Name: 
// Module Name: part_two
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module part_two(
      input reset,
      input clk_in,
      output reg [3:0] redOut,
      output reg [3:0] greenOut,
      output reg [3:0] blueOut,
      output hSync,
      output vSync 
    );
endmodule
